`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 02/06/2021 09:11:04 PM
// Design Name: 
// Module Name: Segment_Seconds
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////




module Segment_Seconds(bcd,seg1);

input [5:0] bcd;
output reg [13:0] seg1;

always @ (bcd)
begin
   case(bcd)
          0: seg1 = 14'b0000001_0000001; // "0"     
          1: seg1 = 14'b0000001_1001111; // "1" 
          2: seg1 = 14'b0000001_0010010; // "2" 
          3: seg1 = 14'b0000001_0000110; // "3" 
          4: seg1 = 14'b0000001_1001100; // "4" 
          5: seg1 = 14'b0000001_0100100; // "5" 
          6: seg1 = 14'b0000001_0100000; // "6" 
          7: seg1 = 14'b0000001_0001111; // "7" 
          8: seg1 = 14'b0000001_0000000; // "8"     
          9: seg1 = 14'b0000001_0000100; // "9"
          
          10: seg1 = 14'b1001111_0000001; // "10"     
          11: seg1 = 14'b1001111_1001111; // "11" 
          12: seg1 = 14'b1001111_0010010; // "12" 
          13: seg1 = 14'b1001111_0000110; // "13" 
          14: seg1 = 14'b1001111_1001100; // "14" 
          15: seg1 = 14'b1001111_0100100; // "15" 
          16: seg1 = 14'b1001111_0100000; // "16" 
          17: seg1 = 14'b1001111_0001111; // "17" 
          18: seg1 = 14'b1001111_0000000; // "18"     
          19: seg1 = 14'b1001111_0000100; // "19"
          
  
          20: seg1 = 14'b0010010_0000001; // "10"     
          21: seg1 = 14'b0010010_1001111; // "11" 
          22: seg1 = 14'b0010010_0010010; // "12" 
          23: seg1 = 14'b0010010_0000110; // "13" 
          24: seg1 = 14'b0010010_1001100; // "14" 
          25: seg1 = 14'b0010010_0100100; // "15" 
          26: seg1 = 14'b0010010_0100000; // "16" 
          27: seg1 = 14'b0010010_0001111; // "17" 
          28: seg1 = 14'b0010010_0000000; // "18"     
          29: seg1 = 14'b0010010_0000100; // "19"


          30: seg1 = 14'b0000110_0000001; // "10"     
          31: seg1 = 14'b0000110_1001111; // "11" 
          32: seg1 = 14'b0000110_0010010; // "12" 
          33: seg1 = 14'b0000110_0000110; // "13" 
          34: seg1 = 14'b0000110_1001100; // "14" 
          35: seg1 = 14'b0000110_0100100; // "15" 
          36: seg1 = 14'b0000110_0100000; // "16" 
          37: seg1 = 14'b0000110_0001111; // "17" 
          38: seg1 = 14'b0000110_0000000; // "18"     
          39: seg1 = 14'b0000110_0000100; // "19"

          40: seg1 = 14'b1001100_0000001; // "10"     
          41: seg1 = 14'b1001100_1001111; // "11" 
          42: seg1 = 14'b1001100_0010010; // "12" 
          43: seg1 = 14'b1001100_0000110; // "13" 
          44: seg1 = 14'b1001100_1001100; // "14" 
          45: seg1 = 14'b1001100_0100100; // "15" 
          46: seg1 = 14'b1001100_0100000; // "16" 
          47: seg1 = 14'b1001100_0001111; // "17" 
          48: seg1 = 14'b1001100_0000000; // "18"     
          49: seg1 = 14'b1001100_0000100; // "19"

          50: seg1 = 14'b0100100_0000001; // "10"     
          51: seg1 = 14'b0100100_1001111; // "11" 
          52: seg1 = 14'b0100100_0010010; // "12" 
          53: seg1 = 14'b0100100_0000110; // "13" 
          54: seg1 = 14'b0100100_1001100; // "14" 
          55: seg1 = 14'b0100100_0100100; // "15" 
          56: seg1 = 14'b0100100_0100000; // "16" 
          57: seg1 = 14'b0100100_0001111; // "17" 
          58: seg1 = 14'b0100100_0000000; // "18"     
          59: seg1 = 14'b0100100_0000100; // "19"
          
          
          
          
          
          
  
          default: seg1 = 14'b0000001_0000001;
    endcase
   
end    

endmodule
